//******************************************************************************
// Time Domain Processing Module
// 
// This module implements the time domain preprocessing for LC3plus encoder,
// including PCM input formatting, pre-emphasis filtering, windowing, and
// overlap-add buffer management.
//
// Features:
// - Multi-channel PCM input processing (1-8 channels)
// - Pre-emphasis filtering with configurable coefficient
// - Hanning window application with 50% overlap
// - Frame segmentation and buffer management
// 
// Author: Audio Codec Design Team
// Date: 2024-06-11
// Version: 1.0
//******************************************************************************

`timescale 1ns/1ps

module time_domain_proc (
    // Clock and reset
    input               clk,
    input               rst_n,
    
    // Control interface
    input               enable,         // Module enable
    input               start,          // Start processing
    output  reg         done,           // Processing complete
    output  reg         error,          // Error flag
    
    // Configuration parameters
    input   [15:0]      frame_length,   // Frame length in samples
    input   [2:0]       channels,       // Number of channels (1-8)
    input   [1:0]       sample_width,   // Sample width: 00=16bit, 01=24bit
    input   [15:0]      preemph_coeff,  // Pre-emphasis coefficient (Q15)
    
    // PCM input data interface
    input   [31:0]      pcm_data,       // PCM input data
    input               pcm_valid,      // PCM data valid
    output  reg         pcm_ready,      // PCM data ready
    
    // Time domain output interface
    output  reg [23:0]  time_data,      // Time domain output (Q23)
    output  reg         time_valid,     // Time domain data valid
    input               time_ready,     // Downstream ready
    
    // Memory interface - Audio buffer
    output  reg [11:0]  mem_addr,       // Memory address
    output  reg [31:0]  mem_wdata,      // Memory write data
    input   [31:0]      mem_rdata,      // Memory read data
    output  reg         mem_wen,        // Memory write enable
    output  reg         mem_ren,        // Memory read enable
    
    // Memory interface - Coefficient ROM
    output  reg [11:0]  coeff_addr,     // Coefficient ROM address
    input   [31:0]      coeff_data,     // Coefficient ROM data
    output  reg         coeff_ren,      // Coefficient ROM read enable
    
    // Debug interface
    output  [31:0]      debug_status
);

    // State machine definitions
    parameter [2:0] IDLE        = 3'b000;
    parameter [2:0] INPUT_PCM   = 3'b001;
    parameter [2:0] PREEMPH     = 3'b010;
    parameter [2:0] WINDOWING   = 3'b011;
    parameter [2:0] OUTPUT      = 3'b100;
    parameter [2:0] ERROR_STATE = 3'b111;
    
    // State registers
    reg [2:0] state, next_state;
    
    // Internal registers
    reg [15:0] sample_count;        // Current sample count
    reg [2:0]  channel_count;       // Current channel
    reg [11:0] buffer_addr;         // Buffer address pointer
    reg [11:0] window_addr;         // Window coefficient address
    reg [31:0] pcm_buffer;          // PCM input buffer
    reg [23:0] preemph_mem;         // Pre-emphasis memory
    reg [31:0] windowed_sample;     // Windowed sample accumulator
    
    // Control flags
    reg input_complete;
    reg preemph_complete;
    reg window_complete;
    reg output_complete;
    
    // Sample format conversion
    reg [23:0] pcm_sample_24bit;
    
    always @(*) begin
        case (sample_width)
            2'b00: pcm_sample_24bit = {{8{pcm_data[15]}}, pcm_data[15:0]};  // 16-bit sign extend
            2'b01: pcm_sample_24bit = pcm_data[23:0];                       // 24-bit direct
            default: pcm_sample_24bit = 24'h000000;
        endcase
    end
    
    // State machine
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
        end else begin
            state <= next_state;
        end
    end
    
    // Next state logic
    always @(*) begin
        case (state)
            IDLE: begin
                if (enable && start) begin
                    next_state = INPUT_PCM;
                end else begin
                    next_state = IDLE;
                end
            end
            
            INPUT_PCM: begin
                if (input_complete) begin
                    next_state = PREEMPH;
                end else if (error) begin
                    next_state = ERROR_STATE;
                end else begin
                    next_state = INPUT_PCM;
                end
            end
            
            PREEMPH: begin
                if (preemph_complete) begin
                    next_state = WINDOWING;
                end else begin
                    next_state = PREEMPH;
                end
            end
            
            WINDOWING: begin
                if (window_complete) begin
                    next_state = OUTPUT;
                end else begin
                    next_state = WINDOWING;
                end
            end
            
            OUTPUT: begin
                if (output_complete) begin
                    next_state = IDLE;
                end else begin
                    next_state = OUTPUT;
                end
            end
            
            ERROR_STATE: begin
                next_state = IDLE;
            end
            
            default: begin
                next_state = IDLE;
            end
        endcase
    end
    
    // PCM input processing
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            sample_count <= 16'h0000;
            channel_count <= 3'b000;
            buffer_addr <= 12'h000;
            input_complete <= 1'b0;
            pcm_ready <= 1'b0;
            mem_wen <= 1'b0;
            mem_addr <= 12'h000;
            mem_wdata <= 32'h00000000;
        end else begin
            case (state)
                IDLE: begin
                    sample_count <= 16'h0000;
                    channel_count <= 3'b000;
                    buffer_addr <= 12'h000;
                    input_complete <= 1'b0;
                    pcm_ready <= enable;
                    mem_wen <= 1'b0;
                end
                
                INPUT_PCM: begin
                    pcm_ready <= 1'b1;
                    
                    if (pcm_valid && pcm_ready) begin
                        // Store PCM sample in buffer
                        mem_addr <= buffer_addr;
                        mem_wdata <= {8'h00, pcm_sample_24bit};
                        mem_wen <= 1'b1;
                        
                        // Update counters
                        if (channel_count == channels) begin
                            channel_count <= 3'b000;
                            sample_count <= sample_count + 1;
                            buffer_addr <= buffer_addr + 1;
                            
                            if (sample_count == frame_length - 1) begin
                                input_complete <= 1'b1;
                                pcm_ready <= 1'b0;
                            end
                        end else begin
                            channel_count <= channel_count + 1;
                            buffer_addr <= buffer_addr + 1;
                        end
                    end else begin
                        mem_wen <= 1'b0;
                    end
                end
                
                default: begin
                    pcm_ready <= 1'b0;
                    mem_wen <= 1'b0;
                end
            endcase
        end
    end
    
    // Pre-emphasis filtering
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            preemph_complete <= 1'b0;
            preemph_mem <= 24'h000000;
            mem_ren <= 1'b0;
        end else begin
            case (state)
                IDLE: begin
                    preemph_complete <= 1'b0;
                    preemph_mem <= 24'h000000;
                    mem_ren <= 1'b0;
                end
                
                PREEMPH: begin
                    // Read sample from buffer
                    mem_addr <= sample_count;
                    mem_ren <= 1'b1;
                    
                    if (mem_ren) begin
                        // Apply pre-emphasis filter: y[n] = x[n] - alpha * x[n-1]
                        // Note: This is a simplified implementation
                        reg [47:0] temp_result;
                        temp_result = mem_rdata[23:0] - ((preemph_coeff * preemph_mem) >>> 15);
                        
                        // Store filtered result back to buffer
                        mem_wdata <= {8'h00, temp_result[23:0]};
                        mem_wen <= 1'b1;
                        
                        // Update pre-emphasis memory
                        preemph_mem <= mem_rdata[23:0];
                        
                        // Update counter
                        sample_count <= sample_count + 1;
                        
                        if (sample_count == frame_length - 1) begin
                            preemph_complete <= 1'b1;
                            mem_ren <= 1'b0;
                            mem_wen <= 1'b0;
                        end
                    end
                end
                
                default: begin
                    mem_ren <= 1'b0;
                end
            endcase
        end
    end
    
    // Windowing operation
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            window_complete <= 1'b0;
            window_addr <= 12'h400;    // Window coefficients start at 0x400
            coeff_ren <= 1'b0;
        end else begin
            case (state)
                IDLE: begin
                    window_complete <= 1'b0;
                    window_addr <= 12'h400;
                    coeff_ren <= 1'b0;
                    sample_count <= 16'h0000;
                end
                
                WINDOWING: begin
                    // Read window coefficient
                    coeff_addr <= window_addr + sample_count;
                    coeff_ren <= 1'b1;
                    
                    // Read sample from buffer
                    mem_addr <= sample_count;
                    mem_ren <= 1'b1;
                    
                    if (coeff_ren && mem_ren) begin
                        // Apply window: windowed = sample * window_coeff
                        reg [55:0] mult_result;
                        mult_result = mem_rdata[23:0] * coeff_data[30:0];  // Q23 * Q31 = Q54
                        windowed_sample <= mult_result[54:31];              // Keep Q23 format
                        
                        // Store windowed result back to buffer
                        mem_wdata <= {8'h00, mult_result[54:31]};
                        mem_wen <= 1'b1;
                        
                        sample_count <= sample_count + 1;
                        
                        if (sample_count == frame_length - 1) begin
                            window_complete <= 1'b1;
                            coeff_ren <= 1'b0;
                            mem_ren <= 1'b0;
                            mem_wen <= 1'b0;
                        end
                    end
                end
                
                default: begin
                    coeff_ren <= 1'b0;
                end
            endcase
        end
    end
    
    // Output data streaming
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            output_complete <= 1'b0;
            time_valid <= 1'b0;
            time_data <= 24'h000000;
        end else begin
            case (state)
                IDLE: begin
                    output_complete <= 1'b0;
                    time_valid <= 1'b0;
                    sample_count <= 16'h0000;
                end
                
                OUTPUT: begin
                    if (time_ready) begin
                        // Read processed sample from buffer
                        mem_addr <= sample_count;
                        mem_ren <= 1'b1;
                        
                        if (mem_ren) begin
                            time_data <= mem_rdata[23:0];
                            time_valid <= 1'b1;
                            
                            sample_count <= sample_count + 1;
                            
                            if (sample_count == frame_length - 1) begin
                                output_complete <= 1'b1;
                                time_valid <= 1'b0;
                                mem_ren <= 1'b0;
                            end
                        end
                    end else begin
                        time_valid <= 1'b0;
                        mem_ren <= 1'b0;
                    end
                end
                
                default: begin
                    time_valid <= 1'b0;
                    mem_ren <= 1'b0;
                end
            endcase
        end
    end
    
    // Status and control signals
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            done <= 1'b0;
            error <= 1'b0;
        end else begin
            case (state)
                IDLE: begin
                    done <= 1'b0;
                    error <= 1'b0;
                end
                
                OUTPUT: begin
                    done <= output_complete;
                end
                
                ERROR_STATE: begin
                    error <= 1'b1;
                end
                
                default: begin
                    done <= 1'b0;
                end
            endcase
        end
    end
    
    // Debug status
    assign debug_status = {
        8'h00,                          // [31:24] Reserved
        state,                          // [23:21] Current state
        channels,                       // [20:18] Channel count
        sample_width,                   // [17:16] Sample width
        sample_count                    // [15:0]  Sample count
    };

endmodule

//******************************************************************************
// Time Domain Processing Module Interface Summary
//
// Clock Domain: Single clock domain (clk)
// Reset: Asynchronous active-low reset (rst_n)
//
// Processing Pipeline:
// 1. PCM Input     - Multi-channel PCM data collection
// 2. Pre-emphasis  - High-frequency boost filtering
// 3. Windowing     - Hanning window application
// 4. Output        - Formatted time domain data output
//
// Memory Usage:
// - Audio Buffer: Stores input PCM and processed samples
// - Coefficient ROM: Window function coefficients (0x400-0x5FF)
//
// Performance:
// - Latency: ~4 * frame_length clock cycles
// - Throughput: 1 sample per clock cycle (output phase)
// - Memory Bandwidth: 2 accesses per sample (read + write)
//
//****************************************************************************** 